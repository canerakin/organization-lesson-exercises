library verilog;
use verilog.vl_types.all;
entity thirty_two_bit_ALU_test_bench is
end thirty_two_bit_ALU_test_bench;
